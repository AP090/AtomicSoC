-- DACpll1.vhd

-- Generated using ACDS version 14.0 200 at 2016.10.25.17:36:38

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity DACpll1 is
	port (
		refclk   : in  std_logic := '0'; --  refclk.clk
		rst      : in  std_logic := '0'; --   reset.reset
		outclk_0 : out std_logic         -- outclk0.clk
	);
end entity DACpll1;

architecture rtl of DACpll1 is
	component DACpll1_0002 is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component DACpll1_0002;

begin

	dacpll1_inst : component DACpll1_0002
		port map (
			refclk   => refclk,   --  refclk.clk
			rst      => rst,      --   reset.reset
			outclk_0 => outclk_0, -- outclk0.clk
			locked   => open      -- (terminated)
		);

end architecture rtl; -- of DACpll1
